-- Joel Brigida
-- CDA 4240C: Digital Design Lab
-- This File Implements the Top Level Wrapper for the Entire Vending Machine.

